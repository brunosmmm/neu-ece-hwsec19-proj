`define SIMON_KEY_WIDTH 128
`define SIMON_MAX_BLOCK_WIDTH 128

`define SIMON_MODE_64_128 1'b0
`define SIMON_MODE_128_128 1'b1

`define SIMON_64_128_WORD_SIZE 32
`define SIMON_64_128_KEY_WORDS (128/`SIMON_64_128_WORD_SIZE)
`define SIMON_128_128_WORD_SIZE 64
`define SIMON_128_128_KEY_WORDS (128/`SIMON_128_128_WORD_SIZE)

`define SIMON_64_128_ROUNDS 44
`define SIMON_128_128_ROUNDS 68

// rotate units
`define ROTATE_MODE_LEFT 0
`define ROTATE_MODE_RIGHT 1
